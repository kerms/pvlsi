library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;        -- for addition & counting
use ieee.numeric_std.all;               -- for type conversions

entity shifter_tb is
end shifter_tb;

architecture shifter_tb_arc of shifter_tb is

begin

end  shifter_tb_arc;